{{NP_NAME}}